library verilog;
use verilog.vl_types.all;
entity DECODER_2x4_vlg_check_tst is
    port(
        o0              : in     vl_logic;
        o1              : in     vl_logic;
        o2              : in     vl_logic;
        o3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DECODER_2x4_vlg_check_tst;
